module xor_wave(
      input wire a,
      input wire b,
      output wire y
);
asiign y=a^b;
endmodule
